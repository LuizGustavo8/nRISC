library verilog;
use verilog.vl_types.all;
entity teste_mdi is
end teste_mdi;
