library verilog;
use verilog.vl_types.all;
entity teste_ULA is
end teste_ULA;
