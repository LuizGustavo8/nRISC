library verilog;
use verilog.vl_types.all;
entity teste_mux is
end teste_mux;
