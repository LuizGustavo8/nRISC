
// Memória de Instrucoes
 module MDI(pc, instruction);  
      input     [7:0]pc;  
      output    [17:0]instruction;  
 
      reg [256:0] mem[17:0];
		
		initial begin
 
//Programa Teste - Calcula a Média dos Valores de um Vetor de Tamanho N
mem[0] = 18'b100000101000001000;
mem[1] = 18'b010000101000000000;
mem[2] = 18'b100000111000001000;
mem[3] = 18'b100000001000000011;
mem[4] = 18'b010111001000000000;
mem[5] = 18'b100000001000000101;
mem[6] = 18'b010111001000000001;
mem[7] = 18'b100000001000000100;
mem[8] = 18'b010111001000000010;
mem[9] = 18'b100000001000000001;
mem[10] = 18'b010111001000000011;
mem[11] = 18'b100000001000000111;
mem[12] = 18'b010111001000000100;
mem[13] = 18'b100000001000000111;
mem[14] = 18'b010111001000000101;
mem[15] = 18'b100000001000001000;
mem[16] = 18'b000110101110000011;
mem[17] = 18'b010000110000000001;
mem[18] = 18'b010111001000000111;
mem[19] = 18'b100000110000000000;
mem[20] = 18'b100000100000000000;
mem[21] = 18'b000100101001000101;
mem[22] = 18'b011001000000011101;
mem[23] = 18'b000111100001000000;
mem[24] = 18'b001001001000000000;
mem[25] = 18'b000110001110000000;
mem[26] = 18'b100100100000000001;
mem[27] = 18'b111000000000010110;
mem[28] = 18'b000110101110000011;
mem[29] = 18'b010000110000000001;

		end
      assign instruction = mem[pc];  
 endmodule 