library verilog;
use verilog.vl_types.all;
entity teste_pc is
end teste_pc;
