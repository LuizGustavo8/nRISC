library verilog;
use verilog.vl_types.all;
entity teste_bdr is
end teste_bdr;
