library verilog;
use verilog.vl_types.all;
entity simulacao is
end simulacao;
