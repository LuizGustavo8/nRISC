library verilog;
use verilog.vl_types.all;
entity teste_cdu is
end teste_cdu;
