library verilog;
use verilog.vl_types.all;
entity teste_mux2 is
end teste_mux2;
