library verilog;
use verilog.vl_types.all;
entity teste_udc is
end teste_udc;
