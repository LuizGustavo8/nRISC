library verilog;
use verilog.vl_types.all;
entity teste_mdd is
end teste_mdd;
